// A test bench for step_one

module step_one_tb();
    wire out;

endmodule
